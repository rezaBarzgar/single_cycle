library verilog;
use verilog.vl_types.all;
entity tbmult is
end tbmult;

library verilog;
use verilog.vl_types.all;
entity Pipeline is
    port(
        clk             : in     vl_logic
    );
end Pipeline;

library verilog;
use verilog.vl_types.all;
entity single_cycle is
    port(
        clk             : in     vl_logic
    );
end single_cycle;

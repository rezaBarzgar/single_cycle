library verilog;
use verilog.vl_types.all;
entity Clk is
    port(
        \out\           : out    vl_logic
    );
end Clk;
